library verilog;
use verilog.vl_types.all;
entity ex03_vlg_vec_tst is
end ex03_vlg_vec_tst;
